`timescale 1ps/100fs
module product_24x24(
	input [23:0] a,
	input [23:0] b,
	output[23:0] [23:0] p 
);
  assign p[0][0] = a[0] & b[0];
assign p[1][0] = a[1] & b[0];
assign p[2][0] = a[2] & b[0];
assign p[3][0] = a[3] & b[0];
assign p[4][0] = a[4] & b[0];
assign p[5][0] = a[5] & b[0];
assign p[6][0] = a[6] & b[0];
assign p[7][0] = a[7] & b[0];
assign p[8][0] = a[8] & b[0];
assign p[9][0] = a[9] & b[0];
assign p[10][0] = a[10] & b[0];
assign p[11][0] = a[11] & b[0];
assign p[12][0] = a[12] & b[0];
assign p[13][0] = a[13] & b[0];
assign p[14][0] = a[14] & b[0];
assign p[15][0] = a[15] & b[0];
assign p[16][0] = a[16] & b[0];
assign p[17][0] = a[17] & b[0];
assign p[18][0] = a[18] & b[0];
assign p[19][0] = a[19] & b[0];
assign p[20][0] = a[20] & b[0];
assign p[21][0] = a[21] & b[0];
assign p[22][0] = a[22] & b[0];
assign p[23][0] = a[23] & b[0];
assign p[0][1] = a[0] & b[1];
assign p[1][1] = a[1] & b[1];
assign p[2][1] = a[2] & b[1];
assign p[3][1] = a[3] & b[1];
assign p[4][1] = a[4] & b[1];
assign p[5][1] = a[5] & b[1];
assign p[6][1] = a[6] & b[1];
assign p[7][1] = a[7] & b[1];
assign p[8][1] = a[8] & b[1];
assign p[9][1] = a[9] & b[1];
assign p[10][1] = a[10] & b[1];
assign p[11][1] = a[11] & b[1];
assign p[12][1] = a[12] & b[1];
assign p[13][1] = a[13] & b[1];
assign p[14][1] = a[14] & b[1];
assign p[15][1] = a[15] & b[1];
assign p[16][1] = a[16] & b[1];
assign p[17][1] = a[17] & b[1];
assign p[18][1] = a[18] & b[1];
assign p[19][1] = a[19] & b[1];
assign p[20][1] = a[20] & b[1];
assign p[21][1] = a[21] & b[1];
assign p[22][1] = a[22] & b[1];
assign p[23][1] = a[23] & b[1];
assign p[0][2] = a[0] & b[2];
assign p[1][2] = a[1] & b[2];
assign p[2][2] = a[2] & b[2];
assign p[3][2] = a[3] & b[2];
assign p[4][2] = a[4] & b[2];
assign p[5][2] = a[5] & b[2];
assign p[6][2] = a[6] & b[2];
assign p[7][2] = a[7] & b[2];
assign p[8][2] = a[8] & b[2];
assign p[9][2] = a[9] & b[2];
assign p[10][2] = a[10] & b[2];
assign p[11][2] = a[11] & b[2];
assign p[12][2] = a[12] & b[2];
assign p[13][2] = a[13] & b[2];
assign p[14][2] = a[14] & b[2];
assign p[15][2] = a[15] & b[2];
assign p[16][2] = a[16] & b[2];
assign p[17][2] = a[17] & b[2];
assign p[18][2] = a[18] & b[2];
assign p[19][2] = a[19] & b[2];
assign p[20][2] = a[20] & b[2];
assign p[21][2] = a[21] & b[2];
assign p[22][2] = a[22] & b[2];
assign p[23][2] = a[23] & b[2];
assign p[0][3] = a[0] & b[3];
assign p[1][3] = a[1] & b[3];
assign p[2][3] = a[2] & b[3];
assign p[3][3] = a[3] & b[3];
assign p[4][3] = a[4] & b[3];
assign p[5][3] = a[5] & b[3];
assign p[6][3] = a[6] & b[3];
assign p[7][3] = a[7] & b[3];
assign p[8][3] = a[8] & b[3];
assign p[9][3] = a[9] & b[3];
assign p[10][3] = a[10] & b[3];
assign p[11][3] = a[11] & b[3];
assign p[12][3] = a[12] & b[3];
assign p[13][3] = a[13] & b[3];
assign p[14][3] = a[14] & b[3];
assign p[15][3] = a[15] & b[3];
assign p[16][3] = a[16] & b[3];
assign p[17][3] = a[17] & b[3];
assign p[18][3] = a[18] & b[3];
assign p[19][3] = a[19] & b[3];
assign p[20][3] = a[20] & b[3];
assign p[21][3] = a[21] & b[3];
assign p[22][3] = a[22] & b[3];
assign p[23][3] = a[23] & b[3];
assign p[0][4] = a[0] & b[4];
assign p[1][4] = a[1] & b[4];
assign p[2][4] = a[2] & b[4];
assign p[3][4] = a[3] & b[4];
assign p[4][4] = a[4] & b[4];
assign p[5][4] = a[5] & b[4];
assign p[6][4] = a[6] & b[4];
assign p[7][4] = a[7] & b[4];
assign p[8][4] = a[8] & b[4];
assign p[9][4] = a[9] & b[4];
assign p[10][4] = a[10] & b[4];
assign p[11][4] = a[11] & b[4];
assign p[12][4] = a[12] & b[4];
assign p[13][4] = a[13] & b[4];
assign p[14][4] = a[14] & b[4];
assign p[15][4] = a[15] & b[4];
assign p[16][4] = a[16] & b[4];
assign p[17][4] = a[17] & b[4];
assign p[18][4] = a[18] & b[4];
assign p[19][4] = a[19] & b[4];
assign p[20][4] = a[20] & b[4];
assign p[21][4] = a[21] & b[4];
assign p[22][4] = a[22] & b[4];
assign p[23][4] = a[23] & b[4];
assign p[0][5] = a[0] & b[5];
assign p[1][5] = a[1] & b[5];
assign p[2][5] = a[2] & b[5];
assign p[3][5] = a[3] & b[5];
assign p[4][5] = a[4] & b[5];
assign p[5][5] = a[5] & b[5];
assign p[6][5] = a[6] & b[5];
assign p[7][5] = a[7] & b[5];
assign p[8][5] = a[8] & b[5];
assign p[9][5] = a[9] & b[5];
assign p[10][5] = a[10] & b[5];
assign p[11][5] = a[11] & b[5];
assign p[12][5] = a[12] & b[5];
assign p[13][5] = a[13] & b[5];
assign p[14][5] = a[14] & b[5];
assign p[15][5] = a[15] & b[5];
assign p[16][5] = a[16] & b[5];
assign p[17][5] = a[17] & b[5];
assign p[18][5] = a[18] & b[5];
assign p[19][5] = a[19] & b[5];
assign p[20][5] = a[20] & b[5];
assign p[21][5] = a[21] & b[5];
assign p[22][5] = a[22] & b[5];
assign p[23][5] = a[23] & b[5];
assign p[0][6] = a[0] & b[6];
assign p[1][6] = a[1] & b[6];
assign p[2][6] = a[2] & b[6];
assign p[3][6] = a[3] & b[6];
assign p[4][6] = a[4] & b[6];
assign p[5][6] = a[5] & b[6];
assign p[6][6] = a[6] & b[6];
assign p[7][6] = a[7] & b[6];
assign p[8][6] = a[8] & b[6];
assign p[9][6] = a[9] & b[6];
assign p[10][6] = a[10] & b[6];
assign p[11][6] = a[11] & b[6];
assign p[12][6] = a[12] & b[6];
assign p[13][6] = a[13] & b[6];
assign p[14][6] = a[14] & b[6];
assign p[15][6] = a[15] & b[6];
assign p[16][6] = a[16] & b[6];
assign p[17][6] = a[17] & b[6];
assign p[18][6] = a[18] & b[6];
assign p[19][6] = a[19] & b[6];
assign p[20][6] = a[20] & b[6];
assign p[21][6] = a[21] & b[6];
assign p[22][6] = a[22] & b[6];
assign p[23][6] = a[23] & b[6];
assign p[0][7] = a[0] & b[7];
assign p[1][7] = a[1] & b[7];
assign p[2][7] = a[2] & b[7];
assign p[3][7] = a[3] & b[7];
assign p[4][7] = a[4] & b[7];
assign p[5][7] = a[5] & b[7];
assign p[6][7] = a[6] & b[7];
assign p[7][7] = a[7] & b[7];
assign p[8][7] = a[8] & b[7];
assign p[9][7] = a[9] & b[7];
assign p[10][7] = a[10] & b[7];
assign p[11][7] = a[11] & b[7];
assign p[12][7] = a[12] & b[7];
assign p[13][7] = a[13] & b[7];
assign p[14][7] = a[14] & b[7];
assign p[15][7] = a[15] & b[7];
assign p[16][7] = a[16] & b[7];
assign p[17][7] = a[17] & b[7];
assign p[18][7] = a[18] & b[7];
assign p[19][7] = a[19] & b[7];
assign p[20][7] = a[20] & b[7];
assign p[21][7] = a[21] & b[7];
assign p[22][7] = a[22] & b[7];
assign p[23][7] = a[23] & b[7];
assign p[0][8] = a[0] & b[8];
assign p[1][8] = a[1] & b[8];
assign p[2][8] = a[2] & b[8];
assign p[3][8] = a[3] & b[8];
assign p[4][8] = a[4] & b[8];
assign p[5][8] = a[5] & b[8];
assign p[6][8] = a[6] & b[8];
assign p[7][8] = a[7] & b[8];
assign p[8][8] = a[8] & b[8];
assign p[9][8] = a[9] & b[8];
assign p[10][8] = a[10] & b[8];
assign p[11][8] = a[11] & b[8];
assign p[12][8] = a[12] & b[8];
assign p[13][8] = a[13] & b[8];
assign p[14][8] = a[14] & b[8];
assign p[15][8] = a[15] & b[8];
assign p[16][8] = a[16] & b[8];
assign p[17][8] = a[17] & b[8];
assign p[18][8] = a[18] & b[8];
assign p[19][8] = a[19] & b[8];
assign p[20][8] = a[20] & b[8];
assign p[21][8] = a[21] & b[8];
assign p[22][8] = a[22] & b[8];
assign p[23][8] = a[23] & b[8];
assign p[0][9] = a[0] & b[9];
assign p[1][9] = a[1] & b[9];
assign p[2][9] = a[2] & b[9];
assign p[3][9] = a[3] & b[9];
assign p[4][9] = a[4] & b[9];
assign p[5][9] = a[5] & b[9];
assign p[6][9] = a[6] & b[9];
assign p[7][9] = a[7] & b[9];
assign p[8][9] = a[8] & b[9];
assign p[9][9] = a[9] & b[9];
assign p[10][9] = a[10] & b[9];
assign p[11][9] = a[11] & b[9];
assign p[12][9] = a[12] & b[9];
assign p[13][9] = a[13] & b[9];
assign p[14][9] = a[14] & b[9];
assign p[15][9] = a[15] & b[9];
assign p[16][9] = a[16] & b[9];
assign p[17][9] = a[17] & b[9];
assign p[18][9] = a[18] & b[9];
assign p[19][9] = a[19] & b[9];
assign p[20][9] = a[20] & b[9];
assign p[21][9] = a[21] & b[9];
assign p[22][9] = a[22] & b[9];
assign p[23][9] = a[23] & b[9];
assign p[0][10] = a[0] & b[10];
assign p[1][10] = a[1] & b[10];
assign p[2][10] = a[2] & b[10];
assign p[3][10] = a[3] & b[10];
assign p[4][10] = a[4] & b[10];
assign p[5][10] = a[5] & b[10];
assign p[6][10] = a[6] & b[10];
assign p[7][10] = a[7] & b[10];
assign p[8][10] = a[8] & b[10];
assign p[9][10] = a[9] & b[10];
assign p[10][10] = a[10] & b[10];
assign p[11][10] = a[11] & b[10];
assign p[12][10] = a[12] & b[10];
assign p[13][10] = a[13] & b[10];
assign p[14][10] = a[14] & b[10];
assign p[15][10] = a[15] & b[10];
assign p[16][10] = a[16] & b[10];
assign p[17][10] = a[17] & b[10];
assign p[18][10] = a[18] & b[10];
assign p[19][10] = a[19] & b[10];
assign p[20][10] = a[20] & b[10];
assign p[21][10] = a[21] & b[10];
assign p[22][10] = a[22] & b[10];
assign p[23][10] = a[23] & b[10];
assign p[0][11] = a[0] & b[11];
assign p[1][11] = a[1] & b[11];
assign p[2][11] = a[2] & b[11];
assign p[3][11] = a[3] & b[11];
assign p[4][11] = a[4] & b[11];
assign p[5][11] = a[5] & b[11];
assign p[6][11] = a[6] & b[11];
assign p[7][11] = a[7] & b[11];
assign p[8][11] = a[8] & b[11];
assign p[9][11] = a[9] & b[11];
assign p[10][11] = a[10] & b[11];
assign p[11][11] = a[11] & b[11];
assign p[12][11] = a[12] & b[11];
assign p[13][11] = a[13] & b[11];
assign p[14][11] = a[14] & b[11];
assign p[15][11] = a[15] & b[11];
assign p[16][11] = a[16] & b[11];
assign p[17][11] = a[17] & b[11];
assign p[18][11] = a[18] & b[11];
assign p[19][11] = a[19] & b[11];
assign p[20][11] = a[20] & b[11];
assign p[21][11] = a[21] & b[11];
assign p[22][11] = a[22] & b[11];
assign p[23][11] = a[23] & b[11];
assign p[0][12] = a[0] & b[12];
assign p[1][12] = a[1] & b[12];
assign p[2][12] = a[2] & b[12];
assign p[3][12] = a[3] & b[12];
assign p[4][12] = a[4] & b[12];
assign p[5][12] = a[5] & b[12];
assign p[6][12] = a[6] & b[12];
assign p[7][12] = a[7] & b[12];
assign p[8][12] = a[8] & b[12];
assign p[9][12] = a[9] & b[12];
assign p[10][12] = a[10] & b[12];
assign p[11][12] = a[11] & b[12];
assign p[12][12] = a[12] & b[12];
assign p[13][12] = a[13] & b[12];
assign p[14][12] = a[14] & b[12];
assign p[15][12] = a[15] & b[12];
assign p[16][12] = a[16] & b[12];
assign p[17][12] = a[17] & b[12];
assign p[18][12] = a[18] & b[12];
assign p[19][12] = a[19] & b[12];
assign p[20][12] = a[20] & b[12];
assign p[21][12] = a[21] & b[12];
assign p[22][12] = a[22] & b[12];
assign p[23][12] = a[23] & b[12];
assign p[0][13] = a[0] & b[13];
assign p[1][13] = a[1] & b[13];
assign p[2][13] = a[2] & b[13];
assign p[3][13] = a[3] & b[13];
assign p[4][13] = a[4] & b[13];
assign p[5][13] = a[5] & b[13];
assign p[6][13] = a[6] & b[13];
assign p[7][13] = a[7] & b[13];
assign p[8][13] = a[8] & b[13];
assign p[9][13] = a[9] & b[13];
assign p[10][13] = a[10] & b[13];
assign p[11][13] = a[11] & b[13];
assign p[12][13] = a[12] & b[13];
assign p[13][13] = a[13] & b[13];
assign p[14][13] = a[14] & b[13];
assign p[15][13] = a[15] & b[13];
assign p[16][13] = a[16] & b[13];
assign p[17][13] = a[17] & b[13];
assign p[18][13] = a[18] & b[13];
assign p[19][13] = a[19] & b[13];
assign p[20][13] = a[20] & b[13];
assign p[21][13] = a[21] & b[13];
assign p[22][13] = a[22] & b[13];
assign p[23][13] = a[23] & b[13];
assign p[0][14] = a[0] & b[14];
assign p[1][14] = a[1] & b[14];
assign p[2][14] = a[2] & b[14];
assign p[3][14] = a[3] & b[14];
assign p[4][14] = a[4] & b[14];
assign p[5][14] = a[5] & b[14];
assign p[6][14] = a[6] & b[14];
assign p[7][14] = a[7] & b[14];
assign p[8][14] = a[8] & b[14];
assign p[9][14] = a[9] & b[14];
assign p[10][14] = a[10] & b[14];
assign p[11][14] = a[11] & b[14];
assign p[12][14] = a[12] & b[14];
assign p[13][14] = a[13] & b[14];
assign p[14][14] = a[14] & b[14];
assign p[15][14] = a[15] & b[14];
assign p[16][14] = a[16] & b[14];
assign p[17][14] = a[17] & b[14];
assign p[18][14] = a[18] & b[14];
assign p[19][14] = a[19] & b[14];
assign p[20][14] = a[20] & b[14];
assign p[21][14] = a[21] & b[14];
assign p[22][14] = a[22] & b[14];
assign p[23][14] = a[23] & b[14];
assign p[0][15] = a[0] & b[15];
assign p[1][15] = a[1] & b[15];
assign p[2][15] = a[2] & b[15];
assign p[3][15] = a[3] & b[15];
assign p[4][15] = a[4] & b[15];
assign p[5][15] = a[5] & b[15];
assign p[6][15] = a[6] & b[15];
assign p[7][15] = a[7] & b[15];
assign p[8][15] = a[8] & b[15];
assign p[9][15] = a[9] & b[15];
assign p[10][15] = a[10] & b[15];
assign p[11][15] = a[11] & b[15];
assign p[12][15] = a[12] & b[15];
assign p[13][15] = a[13] & b[15];
assign p[14][15] = a[14] & b[15];
assign p[15][15] = a[15] & b[15];
assign p[16][15] = a[16] & b[15];
assign p[17][15] = a[17] & b[15];
assign p[18][15] = a[18] & b[15];
assign p[19][15] = a[19] & b[15];
assign p[20][15] = a[20] & b[15];
assign p[21][15] = a[21] & b[15];
assign p[22][15] = a[22] & b[15];
assign p[23][15] = a[23] & b[15];
assign p[0][16] = a[0] & b[16];
assign p[1][16] = a[1] & b[16];
assign p[2][16] = a[2] & b[16];
assign p[3][16] = a[3] & b[16];
assign p[4][16] = a[4] & b[16];
assign p[5][16] = a[5] & b[16];
assign p[6][16] = a[6] & b[16];
assign p[7][16] = a[7] & b[16];
assign p[8][16] = a[8] & b[16];
assign p[9][16] = a[9] & b[16];
assign p[10][16] = a[10] & b[16];
assign p[11][16] = a[11] & b[16];
assign p[12][16] = a[12] & b[16];
assign p[13][16] = a[13] & b[16];
assign p[14][16] = a[14] & b[16];
assign p[15][16] = a[15] & b[16];
assign p[16][16] = a[16] & b[16];
assign p[17][16] = a[17] & b[16];
assign p[18][16] = a[18] & b[16];
assign p[19][16] = a[19] & b[16];
assign p[20][16] = a[20] & b[16];
assign p[21][16] = a[21] & b[16];
assign p[22][16] = a[22] & b[16];
assign p[23][16] = a[23] & b[16];
assign p[0][17] = a[0] & b[17];
assign p[1][17] = a[1] & b[17];
assign p[2][17] = a[2] & b[17];
assign p[3][17] = a[3] & b[17];
assign p[4][17] = a[4] & b[17];
assign p[5][17] = a[5] & b[17];
assign p[6][17] = a[6] & b[17];
assign p[7][17] = a[7] & b[17];
assign p[8][17] = a[8] & b[17];
assign p[9][17] = a[9] & b[17];
assign p[10][17] = a[10] & b[17];
assign p[11][17] = a[11] & b[17];
assign p[12][17] = a[12] & b[17];
assign p[13][17] = a[13] & b[17];
assign p[14][17] = a[14] & b[17];
assign p[15][17] = a[15] & b[17];
assign p[16][17] = a[16] & b[17];
assign p[17][17] = a[17] & b[17];
assign p[18][17] = a[18] & b[17];
assign p[19][17] = a[19] & b[17];
assign p[20][17] = a[20] & b[17];
assign p[21][17] = a[21] & b[17];
assign p[22][17] = a[22] & b[17];
assign p[23][17] = a[23] & b[17];
assign p[0][18] = a[0] & b[18];
assign p[1][18] = a[1] & b[18];
assign p[2][18] = a[2] & b[18];
assign p[3][18] = a[3] & b[18];
assign p[4][18] = a[4] & b[18];
assign p[5][18] = a[5] & b[18];
assign p[6][18] = a[6] & b[18];
assign p[7][18] = a[7] & b[18];
assign p[8][18] = a[8] & b[18];
assign p[9][18] = a[9] & b[18];
assign p[10][18] = a[10] & b[18];
assign p[11][18] = a[11] & b[18];
assign p[12][18] = a[12] & b[18];
assign p[13][18] = a[13] & b[18];
assign p[14][18] = a[14] & b[18];
assign p[15][18] = a[15] & b[18];
assign p[16][18] = a[16] & b[18];
assign p[17][18] = a[17] & b[18];
assign p[18][18] = a[18] & b[18];
assign p[19][18] = a[19] & b[18];
assign p[20][18] = a[20] & b[18];
assign p[21][18] = a[21] & b[18];
assign p[22][18] = a[22] & b[18];
assign p[23][18] = a[23] & b[18];
assign p[0][19] = a[0] & b[19];
assign p[1][19] = a[1] & b[19];
assign p[2][19] = a[2] & b[19];
assign p[3][19] = a[3] & b[19];
assign p[4][19] = a[4] & b[19];
assign p[5][19] = a[5] & b[19];
assign p[6][19] = a[6] & b[19];
assign p[7][19] = a[7] & b[19];
assign p[8][19] = a[8] & b[19];
assign p[9][19] = a[9] & b[19];
assign p[10][19] = a[10] & b[19];
assign p[11][19] = a[11] & b[19];
assign p[12][19] = a[12] & b[19];
assign p[13][19] = a[13] & b[19];
assign p[14][19] = a[14] & b[19];
assign p[15][19] = a[15] & b[19];
assign p[16][19] = a[16] & b[19];
assign p[17][19] = a[17] & b[19];
assign p[18][19] = a[18] & b[19];
assign p[19][19] = a[19] & b[19];
assign p[20][19] = a[20] & b[19];
assign p[21][19] = a[21] & b[19];
assign p[22][19] = a[22] & b[19];
assign p[23][19] = a[23] & b[19];
assign p[0][20] = a[0] & b[20];
assign p[1][20] = a[1] & b[20];
assign p[2][20] = a[2] & b[20];
assign p[3][20] = a[3] & b[20];
assign p[4][20] = a[4] & b[20];
assign p[5][20] = a[5] & b[20];
assign p[6][20] = a[6] & b[20];
assign p[7][20] = a[7] & b[20];
assign p[8][20] = a[8] & b[20];
assign p[9][20] = a[9] & b[20];
assign p[10][20] = a[10] & b[20];
assign p[11][20] = a[11] & b[20];
assign p[12][20] = a[12] & b[20];
assign p[13][20] = a[13] & b[20];
assign p[14][20] = a[14] & b[20];
assign p[15][20] = a[15] & b[20];
assign p[16][20] = a[16] & b[20];
assign p[17][20] = a[17] & b[20];
assign p[18][20] = a[18] & b[20];
assign p[19][20] = a[19] & b[20];
assign p[20][20] = a[20] & b[20];
assign p[21][20] = a[21] & b[20];
assign p[22][20] = a[22] & b[20];
assign p[23][20] = a[23] & b[20];
assign p[0][21] = a[0] & b[21];
assign p[1][21] = a[1] & b[21];
assign p[2][21] = a[2] & b[21];
assign p[3][21] = a[3] & b[21];
assign p[4][21] = a[4] & b[21];
assign p[5][21] = a[5] & b[21];
assign p[6][21] = a[6] & b[21];
assign p[7][21] = a[7] & b[21];
assign p[8][21] = a[8] & b[21];
assign p[9][21] = a[9] & b[21];
assign p[10][21] = a[10] & b[21];
assign p[11][21] = a[11] & b[21];
assign p[12][21] = a[12] & b[21];
assign p[13][21] = a[13] & b[21];
assign p[14][21] = a[14] & b[21];
assign p[15][21] = a[15] & b[21];
assign p[16][21] = a[16] & b[21];
assign p[17][21] = a[17] & b[21];
assign p[18][21] = a[18] & b[21];
assign p[19][21] = a[19] & b[21];
assign p[20][21] = a[20] & b[21];
assign p[21][21] = a[21] & b[21];
assign p[22][21] = a[22] & b[21];
assign p[23][21] = a[23] & b[21];
assign p[0][22] = a[0] & b[22];
assign p[1][22] = a[1] & b[22];
assign p[2][22] = a[2] & b[22];
assign p[3][22] = a[3] & b[22];
assign p[4][22] = a[4] & b[22];
assign p[5][22] = a[5] & b[22];
assign p[6][22] = a[6] & b[22];
assign p[7][22] = a[7] & b[22];
assign p[8][22] = a[8] & b[22];
assign p[9][22] = a[9] & b[22];
assign p[10][22] = a[10] & b[22];
assign p[11][22] = a[11] & b[22];
assign p[12][22] = a[12] & b[22];
assign p[13][22] = a[13] & b[22];
assign p[14][22] = a[14] & b[22];
assign p[15][22] = a[15] & b[22];
assign p[16][22] = a[16] & b[22];
assign p[17][22] = a[17] & b[22];
assign p[18][22] = a[18] & b[22];
assign p[19][22] = a[19] & b[22];
assign p[20][22] = a[20] & b[22];
assign p[21][22] = a[21] & b[22];
assign p[22][22] = a[22] & b[22];
assign p[23][22] = a[23] & b[22];
assign p[0][23] = a[0] & b[23];
assign p[1][23] = a[1] & b[23];
assign p[2][23] = a[2] & b[23];
assign p[3][23] = a[3] & b[23];
assign p[4][23] = a[4] & b[23];
assign p[5][23] = a[5] & b[23];
assign p[6][23] = a[6] & b[23];
assign p[7][23] = a[7] & b[23];
assign p[8][23] = a[8] & b[23];
assign p[9][23] = a[9] & b[23];
assign p[10][23] = a[10] & b[23];
assign p[11][23] = a[11] & b[23];
assign p[12][23] = a[12] & b[23];
assign p[13][23] = a[13] & b[23];
assign p[14][23] = a[14] & b[23];
assign p[15][23] = a[15] & b[23];
assign p[16][23] = a[16] & b[23];
assign p[17][23] = a[17] & b[23];
assign p[18][23] = a[18] & b[23];
assign p[19][23] = a[19] & b[23];
assign p[20][23] = a[20] & b[23];
assign p[21][23] = a[21] & b[23];
assign p[22][23] = a[22] & b[23];
assign p[23][23] = a[23] & b[23];
endmodule
